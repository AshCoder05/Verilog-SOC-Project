// Code your design here
module datapath (
    input wire clk,
    input wire rst,
    
    input wire ld_regs,   
    input wire add_en,    
    input wire shift_en, 
    // Data inputs
    input wire [3:0] multiplier_in,  
    input wire [3:0] multiplicand_in, 
    output wire q0,       
    output wire [7:0] product_out
);
    reg [4:0] A; // 5 bits to handle carry overflow
    reg [3:0] M;
    reg [3:0] Q;

    // LOGIC
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            A <= 0;
            M <= 0;
            Q <= 0;
        end 
        else if (ld_regs) begin
            M <= multiplicand_in;
            Q <= multiplier_in;
            A <= 0; 
        end 
        else begin
            if (add_en) begin
                A <= A + M;
            end
            else if (shift_en) begin
                {A, Q} <= {A, Q} >> 1;
            end
        end
    end

    // CONNECT OUTPUTS
    assign q0 = Q[0];           
    assign product_out = {A[3:0], Q}; 

endmodule

module controller (
    input wire clk, rst, start, q0,
    output reg ld_regs, add_en, shift_en, done
);
    reg [2:0] count;
    reg [2:0] state, next_state;
    
    // States
    parameter S_IDLE=0, S_LOAD=1, S_CHECK=2, S_ADD=3, S_SHIFT=4, S_DONE=5;

    // State Update & Counter
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= S_IDLE;
            count <= 0;
        end else begin
            state <= next_state;
            if (state == S_LOAD) count <= 4;
            else if (state == S_SHIFT) count <= count - 1;
        end
    end

    // Next State Logic
    always @(*) begin
        ld_regs = 0; add_en = 0; shift_en = 0; done = 0;
        next_state = state;

        case (state)
            S_IDLE:  if (start) next_state = S_LOAD;
            S_LOAD:  begin ld_regs=1; next_state = S_CHECK; end
            S_CHECK: if (q0) next_state = S_ADD; else next_state = S_SHIFT;
            S_ADD:   begin add_en=1; next_state = S_SHIFT; end
            S_SHIFT: begin shift_en=1; if(count==1) next_state=S_DONE; else next_state=S_CHECK; end
            S_DONE:  begin done=1; if(!start) next_state = S_IDLE; end
            default: next_state = S_IDLE;
        endcase
    end
endmodule

module sequential_multiplier_top (
    input wire clk, rst, start,
    input wire [3:0] A_in, B_in,
    output wire [7:0] result,
    output wire done
);
    wire ld, add, shift, q0_bit;

    controller Control (
        .clk(clk), .rst(rst), .start(start), .q0(q0_bit),
        .ld_regs(ld), .add_en(add), .shift_en(shift), .done(done)
    );

    datapath Data (
        .clk(clk), .rst(rst), 
        .ld_regs(ld), .add_en(add), .shift_en(shift),
        .multiplier_in(A_in), .multiplicand_in(B_in),
        .q0(q0_bit), .product_out(result)
    );
endmodule
